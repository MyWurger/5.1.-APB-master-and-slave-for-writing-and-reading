// Модуль "СЛЕЙВ"
module slave
#(
  parameter number_in_group_ADDR = 4'h0,  // адрес регистра, где хранится номер студента в группе
  parameter data_ADDR = 4'h4,             // адрес регистра, где хранится дата дд.мм.гг
  parameter surname_ADDR = 4'h8,          // адрес регистра, где хранится первые 4 буквы фамилии
  parameter name_ADDR = 4'hC              // адрес регистра, где хранится первые 4 буквы имени
)          

(
    input wire PWRITE,            // сигнал, выбирающий режим записи или чтения (1 - запись, 0 - чтение)
    input wire PCLK,              // сигнал синхронизации
    input wire PSEL,              // сигнал выбора переферии 
    input wire [31:0] PADDR,      // адрес регистра
    input wire [31:0] PWDATA,     // данные для записи в регистр
    input wire PENABLE,           // сигнал разрешения
    output reg [31:0] PRDATA = 0, // данные, прочитанные из регистра
    output reg PREADY = 0         // сигнал готовности (флаг того, что всё сделано успешно)
);

// Объявляем матрицу OP для хранения регистров
reg [31:0] OP [3:0];              // 0 - number_in_group, 1 - data, 2 - surname, 3 - name

// циклы записи и чтения интерфейса APB для переферийного устройства
// реагирует на входной сигнал и изменение переферийного устройства
always @(posedge PSEL or posedge PCLK) 
begin

    // запись в регистры (выбрано переферийное устройство, сигнал записи, разрешена работа с устройством)
    if (PSEL && PWRITE && PENABLE)
     begin
        // ЗАПИСЬ информации в отведённые ячейки
        case(PADDR)
         number_in_group_ADDR: OP[0] <= PWDATA; // запись по адресу регистра номера человека в группе
         data_ADDR: OP[1] <= PWDATA;            // запись по адресу регистра даты
         surname_ADDR: OP[2] <= PWDATA;         // запись по адресу регистра фамилии
         name_ADDR: OP[3] <= PWDATA;            // запись по адресу регистра имени
        endcase

        PRDATA <=0;                             // записанных данных нет
        PREADY <= 1'd1;                         // устанавливаем флаг заверешения операции
    end

    // ЧТЕНИЕ из регистров (выбрано переферийное устройство, подан сигнал чтения, разрешена работа)
    else if (PSEL && !PWRITE && PENABLE)
    begin
        // чтение информации из отведённых ячеек
        case(PADDR)
         number_in_group_ADDR: PRDATA <= OP[0];  // чтение по адресу номера человека в группе
         data_ADDR: PRDATA <= OP[1];             // чтение по адресу регистра даты
         surname_ADDR: PRDATA <= OP[2];          // чтение по адресу регистра фамилии
         name_ADDR: PRDATA <= OP[3];             // чтение по адресу регистра имени
        endcase

        PREADY <= 1'd1;                          // устанавливаем флаг заверешения операции
    end
   
   // сбрасываем PREADY после выполнения записи или чтения
   if (PREADY)
    begin
      PREADY <= !PREADY;
    end
end

endmodule